magic
tech sky130A
magscale 1 2
timestamp 1640879400
<< obsli1 >>
rect 1104 2159 198812 397681
<< obsm1 >>
rect 1026 2128 198812 397712
<< metal2 >>
rect 16670 399200 16726 400000
rect 49974 399200 50030 400000
rect 83278 399200 83334 400000
rect 116674 399200 116730 400000
rect 149978 399200 150034 400000
rect 183282 399200 183338 400000
rect 7654 0 7710 800
rect 23018 0 23074 800
rect 38382 0 38438 800
rect 53746 0 53802 800
rect 69110 0 69166 800
rect 84566 0 84622 800
rect 99930 0 99986 800
rect 115294 0 115350 800
rect 130658 0 130714 800
rect 146114 0 146170 800
rect 161478 0 161534 800
rect 176842 0 176898 800
rect 192206 0 192262 800
<< obsm2 >>
rect 1030 399144 16614 399265
rect 16782 399144 49918 399265
rect 50086 399144 83222 399265
rect 83390 399144 116618 399265
rect 116786 399144 149922 399265
rect 150090 399144 183226 399265
rect 183394 399144 198058 399265
rect 1030 856 198058 399144
rect 1030 575 7598 856
rect 7766 575 22962 856
rect 23130 575 38326 856
rect 38494 575 53690 856
rect 53858 575 69054 856
rect 69222 575 84510 856
rect 84678 575 99874 856
rect 100042 575 115238 856
rect 115406 575 130602 856
rect 130770 575 146058 856
rect 146226 575 161422 856
rect 161590 575 176786 856
rect 176954 575 192150 856
rect 192318 575 198058 856
<< metal3 >>
rect 0 399168 800 399288
rect 0 397808 800 397928
rect 0 396448 800 396568
rect 0 395224 800 395344
rect 0 393864 800 393984
rect 0 392504 800 392624
rect 0 391280 800 391400
rect 0 389920 800 390040
rect 0 388560 800 388680
rect 0 387336 800 387456
rect 0 385976 800 386096
rect 0 384616 800 384736
rect 0 383392 800 383512
rect 0 382032 800 382152
rect 0 380672 800 380792
rect 199200 379856 200000 379976
rect 0 379448 800 379568
rect 0 378088 800 378208
rect 0 376728 800 376848
rect 0 375504 800 375624
rect 0 374144 800 374264
rect 0 372784 800 372904
rect 0 371560 800 371680
rect 0 370200 800 370320
rect 0 368840 800 368960
rect 0 367616 800 367736
rect 0 366256 800 366376
rect 0 364896 800 365016
rect 0 363672 800 363792
rect 0 362312 800 362432
rect 0 360952 800 361072
rect 0 359728 800 359848
rect 0 358368 800 358488
rect 0 357008 800 357128
rect 0 355784 800 355904
rect 0 354424 800 354544
rect 0 353064 800 353184
rect 0 351840 800 351960
rect 0 350480 800 350600
rect 0 349120 800 349240
rect 0 347896 800 348016
rect 0 346536 800 346656
rect 0 345176 800 345296
rect 0 343952 800 344072
rect 0 342592 800 342712
rect 0 341232 800 341352
rect 0 339872 800 339992
rect 199200 339872 200000 339992
rect 0 338648 800 338768
rect 0 337288 800 337408
rect 0 335928 800 336048
rect 0 334704 800 334824
rect 0 333344 800 333464
rect 0 331984 800 332104
rect 0 330760 800 330880
rect 0 329400 800 329520
rect 0 328040 800 328160
rect 0 326816 800 326936
rect 0 325456 800 325576
rect 0 324096 800 324216
rect 0 322872 800 322992
rect 0 321512 800 321632
rect 0 320152 800 320272
rect 0 318928 800 319048
rect 0 317568 800 317688
rect 0 316208 800 316328
rect 0 314984 800 315104
rect 0 313624 800 313744
rect 0 312264 800 312384
rect 0 311040 800 311160
rect 0 309680 800 309800
rect 0 308320 800 308440
rect 0 307096 800 307216
rect 0 305736 800 305856
rect 0 304376 800 304496
rect 0 303152 800 303272
rect 0 301792 800 301912
rect 0 300432 800 300552
rect 199200 299888 200000 300008
rect 0 299208 800 299328
rect 0 297848 800 297968
rect 0 296488 800 296608
rect 0 295264 800 295384
rect 0 293904 800 294024
rect 0 292544 800 292664
rect 0 291320 800 291440
rect 0 289960 800 290080
rect 0 288600 800 288720
rect 0 287376 800 287496
rect 0 286016 800 286136
rect 0 284656 800 284776
rect 0 283296 800 283416
rect 0 282072 800 282192
rect 0 280712 800 280832
rect 0 279352 800 279472
rect 0 278128 800 278248
rect 0 276768 800 276888
rect 0 275408 800 275528
rect 0 274184 800 274304
rect 0 272824 800 272944
rect 0 271464 800 271584
rect 0 270240 800 270360
rect 0 268880 800 269000
rect 0 267520 800 267640
rect 0 266296 800 266416
rect 0 264936 800 265056
rect 0 263576 800 263696
rect 0 262352 800 262472
rect 0 260992 800 261112
rect 199200 259904 200000 260024
rect 0 259632 800 259752
rect 0 258408 800 258528
rect 0 257048 800 257168
rect 0 255688 800 255808
rect 0 254464 800 254584
rect 0 253104 800 253224
rect 0 251744 800 251864
rect 0 250520 800 250640
rect 0 249160 800 249280
rect 0 247800 800 247920
rect 0 246576 800 246696
rect 0 245216 800 245336
rect 0 243856 800 243976
rect 0 242632 800 242752
rect 0 241272 800 241392
rect 0 239912 800 240032
rect 0 238688 800 238808
rect 0 237328 800 237448
rect 0 235968 800 236088
rect 0 234744 800 234864
rect 0 233384 800 233504
rect 0 232024 800 232144
rect 0 230800 800 230920
rect 0 229440 800 229560
rect 0 228080 800 228200
rect 0 226720 800 226840
rect 0 225496 800 225616
rect 0 224136 800 224256
rect 0 222776 800 222896
rect 0 221552 800 221672
rect 0 220192 800 220312
rect 199200 219920 200000 220040
rect 0 218832 800 218952
rect 0 217608 800 217728
rect 0 216248 800 216368
rect 0 214888 800 215008
rect 0 213664 800 213784
rect 0 212304 800 212424
rect 0 210944 800 211064
rect 0 209720 800 209840
rect 0 208360 800 208480
rect 0 207000 800 207120
rect 0 205776 800 205896
rect 0 204416 800 204536
rect 0 203056 800 203176
rect 0 201832 800 201952
rect 0 200472 800 200592
rect 0 199112 800 199232
rect 0 197888 800 198008
rect 0 196528 800 196648
rect 0 195168 800 195288
rect 0 193944 800 194064
rect 0 192584 800 192704
rect 0 191224 800 191344
rect 0 190000 800 190120
rect 0 188640 800 188760
rect 0 187280 800 187400
rect 0 186056 800 186176
rect 0 184696 800 184816
rect 0 183336 800 183456
rect 0 182112 800 182232
rect 0 180752 800 180872
rect 199200 179936 200000 180056
rect 0 179392 800 179512
rect 0 178168 800 178288
rect 0 176808 800 176928
rect 0 175448 800 175568
rect 0 174224 800 174344
rect 0 172864 800 172984
rect 0 171504 800 171624
rect 0 170144 800 170264
rect 0 168920 800 169040
rect 0 167560 800 167680
rect 0 166200 800 166320
rect 0 164976 800 165096
rect 0 163616 800 163736
rect 0 162256 800 162376
rect 0 161032 800 161152
rect 0 159672 800 159792
rect 0 158312 800 158432
rect 0 157088 800 157208
rect 0 155728 800 155848
rect 0 154368 800 154488
rect 0 153144 800 153264
rect 0 151784 800 151904
rect 0 150424 800 150544
rect 0 149200 800 149320
rect 0 147840 800 147960
rect 0 146480 800 146600
rect 0 145256 800 145376
rect 0 143896 800 144016
rect 0 142536 800 142656
rect 0 141312 800 141432
rect 0 139952 800 140072
rect 199200 139952 200000 140072
rect 0 138592 800 138712
rect 0 137368 800 137488
rect 0 136008 800 136128
rect 0 134648 800 134768
rect 0 133424 800 133544
rect 0 132064 800 132184
rect 0 130704 800 130824
rect 0 129480 800 129600
rect 0 128120 800 128240
rect 0 126760 800 126880
rect 0 125536 800 125656
rect 0 124176 800 124296
rect 0 122816 800 122936
rect 0 121592 800 121712
rect 0 120232 800 120352
rect 0 118872 800 118992
rect 0 117648 800 117768
rect 0 116288 800 116408
rect 0 114928 800 115048
rect 0 113568 800 113688
rect 0 112344 800 112464
rect 0 110984 800 111104
rect 0 109624 800 109744
rect 0 108400 800 108520
rect 0 107040 800 107160
rect 0 105680 800 105800
rect 0 104456 800 104576
rect 0 103096 800 103216
rect 0 101736 800 101856
rect 0 100512 800 100632
rect 199200 99968 200000 100088
rect 0 99152 800 99272
rect 0 97792 800 97912
rect 0 96568 800 96688
rect 0 95208 800 95328
rect 0 93848 800 93968
rect 0 92624 800 92744
rect 0 91264 800 91384
rect 0 89904 800 90024
rect 0 88680 800 88800
rect 0 87320 800 87440
rect 0 85960 800 86080
rect 0 84736 800 84856
rect 0 83376 800 83496
rect 0 82016 800 82136
rect 0 80792 800 80912
rect 0 79432 800 79552
rect 0 78072 800 78192
rect 0 76848 800 76968
rect 0 75488 800 75608
rect 0 74128 800 74248
rect 0 72904 800 73024
rect 0 71544 800 71664
rect 0 70184 800 70304
rect 0 68960 800 69080
rect 0 67600 800 67720
rect 0 66240 800 66360
rect 0 65016 800 65136
rect 0 63656 800 63776
rect 0 62296 800 62416
rect 0 61072 800 61192
rect 199200 59984 200000 60104
rect 0 59712 800 59832
rect 0 58352 800 58472
rect 0 56992 800 57112
rect 0 55768 800 55888
rect 0 54408 800 54528
rect 0 53048 800 53168
rect 0 51824 800 51944
rect 0 50464 800 50584
rect 0 49104 800 49224
rect 0 47880 800 48000
rect 0 46520 800 46640
rect 0 45160 800 45280
rect 0 43936 800 44056
rect 0 42576 800 42696
rect 0 41216 800 41336
rect 0 39992 800 40112
rect 0 38632 800 38752
rect 0 37272 800 37392
rect 0 36048 800 36168
rect 0 34688 800 34808
rect 0 33328 800 33448
rect 0 32104 800 32224
rect 0 30744 800 30864
rect 0 29384 800 29504
rect 0 28160 800 28280
rect 0 26800 800 26920
rect 0 25440 800 25560
rect 0 24216 800 24336
rect 0 22856 800 22976
rect 0 21496 800 21616
rect 0 20272 800 20392
rect 199200 20000 200000 20120
rect 0 18912 800 19032
rect 0 17552 800 17672
rect 0 16328 800 16448
rect 0 14968 800 15088
rect 0 13608 800 13728
rect 0 12384 800 12504
rect 0 11024 800 11144
rect 0 9664 800 9784
rect 0 8440 800 8560
rect 0 7080 800 7200
rect 0 5720 800 5840
rect 0 4496 800 4616
rect 0 3136 800 3256
rect 0 1776 800 1896
rect 0 552 800 672
<< obsm3 >>
rect 880 399088 199200 399261
rect 800 398008 199200 399088
rect 880 397728 199200 398008
rect 800 396648 199200 397728
rect 880 396368 199200 396648
rect 800 395424 199200 396368
rect 880 395144 199200 395424
rect 800 394064 199200 395144
rect 880 393784 199200 394064
rect 800 392704 199200 393784
rect 880 392424 199200 392704
rect 800 391480 199200 392424
rect 880 391200 199200 391480
rect 800 390120 199200 391200
rect 880 389840 199200 390120
rect 800 388760 199200 389840
rect 880 388480 199200 388760
rect 800 387536 199200 388480
rect 880 387256 199200 387536
rect 800 386176 199200 387256
rect 880 385896 199200 386176
rect 800 384816 199200 385896
rect 880 384536 199200 384816
rect 800 383592 199200 384536
rect 880 383312 199200 383592
rect 800 382232 199200 383312
rect 880 381952 199200 382232
rect 800 380872 199200 381952
rect 880 380592 199200 380872
rect 800 380056 199200 380592
rect 800 379776 199120 380056
rect 800 379648 199200 379776
rect 880 379368 199200 379648
rect 800 378288 199200 379368
rect 880 378008 199200 378288
rect 800 376928 199200 378008
rect 880 376648 199200 376928
rect 800 375704 199200 376648
rect 880 375424 199200 375704
rect 800 374344 199200 375424
rect 880 374064 199200 374344
rect 800 372984 199200 374064
rect 880 372704 199200 372984
rect 800 371760 199200 372704
rect 880 371480 199200 371760
rect 800 370400 199200 371480
rect 880 370120 199200 370400
rect 800 369040 199200 370120
rect 880 368760 199200 369040
rect 800 367816 199200 368760
rect 880 367536 199200 367816
rect 800 366456 199200 367536
rect 880 366176 199200 366456
rect 800 365096 199200 366176
rect 880 364816 199200 365096
rect 800 363872 199200 364816
rect 880 363592 199200 363872
rect 800 362512 199200 363592
rect 880 362232 199200 362512
rect 800 361152 199200 362232
rect 880 360872 199200 361152
rect 800 359928 199200 360872
rect 880 359648 199200 359928
rect 800 358568 199200 359648
rect 880 358288 199200 358568
rect 800 357208 199200 358288
rect 880 356928 199200 357208
rect 800 355984 199200 356928
rect 880 355704 199200 355984
rect 800 354624 199200 355704
rect 880 354344 199200 354624
rect 800 353264 199200 354344
rect 880 352984 199200 353264
rect 800 352040 199200 352984
rect 880 351760 199200 352040
rect 800 350680 199200 351760
rect 880 350400 199200 350680
rect 800 349320 199200 350400
rect 880 349040 199200 349320
rect 800 348096 199200 349040
rect 880 347816 199200 348096
rect 800 346736 199200 347816
rect 880 346456 199200 346736
rect 800 345376 199200 346456
rect 880 345096 199200 345376
rect 800 344152 199200 345096
rect 880 343872 199200 344152
rect 800 342792 199200 343872
rect 880 342512 199200 342792
rect 800 341432 199200 342512
rect 880 341152 199200 341432
rect 800 340072 199200 341152
rect 880 339792 199120 340072
rect 800 338848 199200 339792
rect 880 338568 199200 338848
rect 800 337488 199200 338568
rect 880 337208 199200 337488
rect 800 336128 199200 337208
rect 880 335848 199200 336128
rect 800 334904 199200 335848
rect 880 334624 199200 334904
rect 800 333544 199200 334624
rect 880 333264 199200 333544
rect 800 332184 199200 333264
rect 880 331904 199200 332184
rect 800 330960 199200 331904
rect 880 330680 199200 330960
rect 800 329600 199200 330680
rect 880 329320 199200 329600
rect 800 328240 199200 329320
rect 880 327960 199200 328240
rect 800 327016 199200 327960
rect 880 326736 199200 327016
rect 800 325656 199200 326736
rect 880 325376 199200 325656
rect 800 324296 199200 325376
rect 880 324016 199200 324296
rect 800 323072 199200 324016
rect 880 322792 199200 323072
rect 800 321712 199200 322792
rect 880 321432 199200 321712
rect 800 320352 199200 321432
rect 880 320072 199200 320352
rect 800 319128 199200 320072
rect 880 318848 199200 319128
rect 800 317768 199200 318848
rect 880 317488 199200 317768
rect 800 316408 199200 317488
rect 880 316128 199200 316408
rect 800 315184 199200 316128
rect 880 314904 199200 315184
rect 800 313824 199200 314904
rect 880 313544 199200 313824
rect 800 312464 199200 313544
rect 880 312184 199200 312464
rect 800 311240 199200 312184
rect 880 310960 199200 311240
rect 800 309880 199200 310960
rect 880 309600 199200 309880
rect 800 308520 199200 309600
rect 880 308240 199200 308520
rect 800 307296 199200 308240
rect 880 307016 199200 307296
rect 800 305936 199200 307016
rect 880 305656 199200 305936
rect 800 304576 199200 305656
rect 880 304296 199200 304576
rect 800 303352 199200 304296
rect 880 303072 199200 303352
rect 800 301992 199200 303072
rect 880 301712 199200 301992
rect 800 300632 199200 301712
rect 880 300352 199200 300632
rect 800 300088 199200 300352
rect 800 299808 199120 300088
rect 800 299408 199200 299808
rect 880 299128 199200 299408
rect 800 298048 199200 299128
rect 880 297768 199200 298048
rect 800 296688 199200 297768
rect 880 296408 199200 296688
rect 800 295464 199200 296408
rect 880 295184 199200 295464
rect 800 294104 199200 295184
rect 880 293824 199200 294104
rect 800 292744 199200 293824
rect 880 292464 199200 292744
rect 800 291520 199200 292464
rect 880 291240 199200 291520
rect 800 290160 199200 291240
rect 880 289880 199200 290160
rect 800 288800 199200 289880
rect 880 288520 199200 288800
rect 800 287576 199200 288520
rect 880 287296 199200 287576
rect 800 286216 199200 287296
rect 880 285936 199200 286216
rect 800 284856 199200 285936
rect 880 284576 199200 284856
rect 800 283496 199200 284576
rect 880 283216 199200 283496
rect 800 282272 199200 283216
rect 880 281992 199200 282272
rect 800 280912 199200 281992
rect 880 280632 199200 280912
rect 800 279552 199200 280632
rect 880 279272 199200 279552
rect 800 278328 199200 279272
rect 880 278048 199200 278328
rect 800 276968 199200 278048
rect 880 276688 199200 276968
rect 800 275608 199200 276688
rect 880 275328 199200 275608
rect 800 274384 199200 275328
rect 880 274104 199200 274384
rect 800 273024 199200 274104
rect 880 272744 199200 273024
rect 800 271664 199200 272744
rect 880 271384 199200 271664
rect 800 270440 199200 271384
rect 880 270160 199200 270440
rect 800 269080 199200 270160
rect 880 268800 199200 269080
rect 800 267720 199200 268800
rect 880 267440 199200 267720
rect 800 266496 199200 267440
rect 880 266216 199200 266496
rect 800 265136 199200 266216
rect 880 264856 199200 265136
rect 800 263776 199200 264856
rect 880 263496 199200 263776
rect 800 262552 199200 263496
rect 880 262272 199200 262552
rect 800 261192 199200 262272
rect 880 260912 199200 261192
rect 800 260104 199200 260912
rect 800 259832 199120 260104
rect 880 259824 199120 259832
rect 880 259552 199200 259824
rect 800 258608 199200 259552
rect 880 258328 199200 258608
rect 800 257248 199200 258328
rect 880 256968 199200 257248
rect 800 255888 199200 256968
rect 880 255608 199200 255888
rect 800 254664 199200 255608
rect 880 254384 199200 254664
rect 800 253304 199200 254384
rect 880 253024 199200 253304
rect 800 251944 199200 253024
rect 880 251664 199200 251944
rect 800 250720 199200 251664
rect 880 250440 199200 250720
rect 800 249360 199200 250440
rect 880 249080 199200 249360
rect 800 248000 199200 249080
rect 880 247720 199200 248000
rect 800 246776 199200 247720
rect 880 246496 199200 246776
rect 800 245416 199200 246496
rect 880 245136 199200 245416
rect 800 244056 199200 245136
rect 880 243776 199200 244056
rect 800 242832 199200 243776
rect 880 242552 199200 242832
rect 800 241472 199200 242552
rect 880 241192 199200 241472
rect 800 240112 199200 241192
rect 880 239832 199200 240112
rect 800 238888 199200 239832
rect 880 238608 199200 238888
rect 800 237528 199200 238608
rect 880 237248 199200 237528
rect 800 236168 199200 237248
rect 880 235888 199200 236168
rect 800 234944 199200 235888
rect 880 234664 199200 234944
rect 800 233584 199200 234664
rect 880 233304 199200 233584
rect 800 232224 199200 233304
rect 880 231944 199200 232224
rect 800 231000 199200 231944
rect 880 230720 199200 231000
rect 800 229640 199200 230720
rect 880 229360 199200 229640
rect 800 228280 199200 229360
rect 880 228000 199200 228280
rect 800 226920 199200 228000
rect 880 226640 199200 226920
rect 800 225696 199200 226640
rect 880 225416 199200 225696
rect 800 224336 199200 225416
rect 880 224056 199200 224336
rect 800 222976 199200 224056
rect 880 222696 199200 222976
rect 800 221752 199200 222696
rect 880 221472 199200 221752
rect 800 220392 199200 221472
rect 880 220120 199200 220392
rect 880 220112 199120 220120
rect 800 219840 199120 220112
rect 800 219032 199200 219840
rect 880 218752 199200 219032
rect 800 217808 199200 218752
rect 880 217528 199200 217808
rect 800 216448 199200 217528
rect 880 216168 199200 216448
rect 800 215088 199200 216168
rect 880 214808 199200 215088
rect 800 213864 199200 214808
rect 880 213584 199200 213864
rect 800 212504 199200 213584
rect 880 212224 199200 212504
rect 800 211144 199200 212224
rect 880 210864 199200 211144
rect 800 209920 199200 210864
rect 880 209640 199200 209920
rect 800 208560 199200 209640
rect 880 208280 199200 208560
rect 800 207200 199200 208280
rect 880 206920 199200 207200
rect 800 205976 199200 206920
rect 880 205696 199200 205976
rect 800 204616 199200 205696
rect 880 204336 199200 204616
rect 800 203256 199200 204336
rect 880 202976 199200 203256
rect 800 202032 199200 202976
rect 880 201752 199200 202032
rect 800 200672 199200 201752
rect 880 200392 199200 200672
rect 800 199312 199200 200392
rect 880 199032 199200 199312
rect 800 198088 199200 199032
rect 880 197808 199200 198088
rect 800 196728 199200 197808
rect 880 196448 199200 196728
rect 800 195368 199200 196448
rect 880 195088 199200 195368
rect 800 194144 199200 195088
rect 880 193864 199200 194144
rect 800 192784 199200 193864
rect 880 192504 199200 192784
rect 800 191424 199200 192504
rect 880 191144 199200 191424
rect 800 190200 199200 191144
rect 880 189920 199200 190200
rect 800 188840 199200 189920
rect 880 188560 199200 188840
rect 800 187480 199200 188560
rect 880 187200 199200 187480
rect 800 186256 199200 187200
rect 880 185976 199200 186256
rect 800 184896 199200 185976
rect 880 184616 199200 184896
rect 800 183536 199200 184616
rect 880 183256 199200 183536
rect 800 182312 199200 183256
rect 880 182032 199200 182312
rect 800 180952 199200 182032
rect 880 180672 199200 180952
rect 800 180136 199200 180672
rect 800 179856 199120 180136
rect 800 179592 199200 179856
rect 880 179312 199200 179592
rect 800 178368 199200 179312
rect 880 178088 199200 178368
rect 800 177008 199200 178088
rect 880 176728 199200 177008
rect 800 175648 199200 176728
rect 880 175368 199200 175648
rect 800 174424 199200 175368
rect 880 174144 199200 174424
rect 800 173064 199200 174144
rect 880 172784 199200 173064
rect 800 171704 199200 172784
rect 880 171424 199200 171704
rect 800 170344 199200 171424
rect 880 170064 199200 170344
rect 800 169120 199200 170064
rect 880 168840 199200 169120
rect 800 167760 199200 168840
rect 880 167480 199200 167760
rect 800 166400 199200 167480
rect 880 166120 199200 166400
rect 800 165176 199200 166120
rect 880 164896 199200 165176
rect 800 163816 199200 164896
rect 880 163536 199200 163816
rect 800 162456 199200 163536
rect 880 162176 199200 162456
rect 800 161232 199200 162176
rect 880 160952 199200 161232
rect 800 159872 199200 160952
rect 880 159592 199200 159872
rect 800 158512 199200 159592
rect 880 158232 199200 158512
rect 800 157288 199200 158232
rect 880 157008 199200 157288
rect 800 155928 199200 157008
rect 880 155648 199200 155928
rect 800 154568 199200 155648
rect 880 154288 199200 154568
rect 800 153344 199200 154288
rect 880 153064 199200 153344
rect 800 151984 199200 153064
rect 880 151704 199200 151984
rect 800 150624 199200 151704
rect 880 150344 199200 150624
rect 800 149400 199200 150344
rect 880 149120 199200 149400
rect 800 148040 199200 149120
rect 880 147760 199200 148040
rect 800 146680 199200 147760
rect 880 146400 199200 146680
rect 800 145456 199200 146400
rect 880 145176 199200 145456
rect 800 144096 199200 145176
rect 880 143816 199200 144096
rect 800 142736 199200 143816
rect 880 142456 199200 142736
rect 800 141512 199200 142456
rect 880 141232 199200 141512
rect 800 140152 199200 141232
rect 880 139872 199120 140152
rect 800 138792 199200 139872
rect 880 138512 199200 138792
rect 800 137568 199200 138512
rect 880 137288 199200 137568
rect 800 136208 199200 137288
rect 880 135928 199200 136208
rect 800 134848 199200 135928
rect 880 134568 199200 134848
rect 800 133624 199200 134568
rect 880 133344 199200 133624
rect 800 132264 199200 133344
rect 880 131984 199200 132264
rect 800 130904 199200 131984
rect 880 130624 199200 130904
rect 800 129680 199200 130624
rect 880 129400 199200 129680
rect 800 128320 199200 129400
rect 880 128040 199200 128320
rect 800 126960 199200 128040
rect 880 126680 199200 126960
rect 800 125736 199200 126680
rect 880 125456 199200 125736
rect 800 124376 199200 125456
rect 880 124096 199200 124376
rect 800 123016 199200 124096
rect 880 122736 199200 123016
rect 800 121792 199200 122736
rect 880 121512 199200 121792
rect 800 120432 199200 121512
rect 880 120152 199200 120432
rect 800 119072 199200 120152
rect 880 118792 199200 119072
rect 800 117848 199200 118792
rect 880 117568 199200 117848
rect 800 116488 199200 117568
rect 880 116208 199200 116488
rect 800 115128 199200 116208
rect 880 114848 199200 115128
rect 800 113768 199200 114848
rect 880 113488 199200 113768
rect 800 112544 199200 113488
rect 880 112264 199200 112544
rect 800 111184 199200 112264
rect 880 110904 199200 111184
rect 800 109824 199200 110904
rect 880 109544 199200 109824
rect 800 108600 199200 109544
rect 880 108320 199200 108600
rect 800 107240 199200 108320
rect 880 106960 199200 107240
rect 800 105880 199200 106960
rect 880 105600 199200 105880
rect 800 104656 199200 105600
rect 880 104376 199200 104656
rect 800 103296 199200 104376
rect 880 103016 199200 103296
rect 800 101936 199200 103016
rect 880 101656 199200 101936
rect 800 100712 199200 101656
rect 880 100432 199200 100712
rect 800 100168 199200 100432
rect 800 99888 199120 100168
rect 800 99352 199200 99888
rect 880 99072 199200 99352
rect 800 97992 199200 99072
rect 880 97712 199200 97992
rect 800 96768 199200 97712
rect 880 96488 199200 96768
rect 800 95408 199200 96488
rect 880 95128 199200 95408
rect 800 94048 199200 95128
rect 880 93768 199200 94048
rect 800 92824 199200 93768
rect 880 92544 199200 92824
rect 800 91464 199200 92544
rect 880 91184 199200 91464
rect 800 90104 199200 91184
rect 880 89824 199200 90104
rect 800 88880 199200 89824
rect 880 88600 199200 88880
rect 800 87520 199200 88600
rect 880 87240 199200 87520
rect 800 86160 199200 87240
rect 880 85880 199200 86160
rect 800 84936 199200 85880
rect 880 84656 199200 84936
rect 800 83576 199200 84656
rect 880 83296 199200 83576
rect 800 82216 199200 83296
rect 880 81936 199200 82216
rect 800 80992 199200 81936
rect 880 80712 199200 80992
rect 800 79632 199200 80712
rect 880 79352 199200 79632
rect 800 78272 199200 79352
rect 880 77992 199200 78272
rect 800 77048 199200 77992
rect 880 76768 199200 77048
rect 800 75688 199200 76768
rect 880 75408 199200 75688
rect 800 74328 199200 75408
rect 880 74048 199200 74328
rect 800 73104 199200 74048
rect 880 72824 199200 73104
rect 800 71744 199200 72824
rect 880 71464 199200 71744
rect 800 70384 199200 71464
rect 880 70104 199200 70384
rect 800 69160 199200 70104
rect 880 68880 199200 69160
rect 800 67800 199200 68880
rect 880 67520 199200 67800
rect 800 66440 199200 67520
rect 880 66160 199200 66440
rect 800 65216 199200 66160
rect 880 64936 199200 65216
rect 800 63856 199200 64936
rect 880 63576 199200 63856
rect 800 62496 199200 63576
rect 880 62216 199200 62496
rect 800 61272 199200 62216
rect 880 60992 199200 61272
rect 800 60184 199200 60992
rect 800 59912 199120 60184
rect 880 59904 199120 59912
rect 880 59632 199200 59904
rect 800 58552 199200 59632
rect 880 58272 199200 58552
rect 800 57192 199200 58272
rect 880 56912 199200 57192
rect 800 55968 199200 56912
rect 880 55688 199200 55968
rect 800 54608 199200 55688
rect 880 54328 199200 54608
rect 800 53248 199200 54328
rect 880 52968 199200 53248
rect 800 52024 199200 52968
rect 880 51744 199200 52024
rect 800 50664 199200 51744
rect 880 50384 199200 50664
rect 800 49304 199200 50384
rect 880 49024 199200 49304
rect 800 48080 199200 49024
rect 880 47800 199200 48080
rect 800 46720 199200 47800
rect 880 46440 199200 46720
rect 800 45360 199200 46440
rect 880 45080 199200 45360
rect 800 44136 199200 45080
rect 880 43856 199200 44136
rect 800 42776 199200 43856
rect 880 42496 199200 42776
rect 800 41416 199200 42496
rect 880 41136 199200 41416
rect 800 40192 199200 41136
rect 880 39912 199200 40192
rect 800 38832 199200 39912
rect 880 38552 199200 38832
rect 800 37472 199200 38552
rect 880 37192 199200 37472
rect 800 36248 199200 37192
rect 880 35968 199200 36248
rect 800 34888 199200 35968
rect 880 34608 199200 34888
rect 800 33528 199200 34608
rect 880 33248 199200 33528
rect 800 32304 199200 33248
rect 880 32024 199200 32304
rect 800 30944 199200 32024
rect 880 30664 199200 30944
rect 800 29584 199200 30664
rect 880 29304 199200 29584
rect 800 28360 199200 29304
rect 880 28080 199200 28360
rect 800 27000 199200 28080
rect 880 26720 199200 27000
rect 800 25640 199200 26720
rect 880 25360 199200 25640
rect 800 24416 199200 25360
rect 880 24136 199200 24416
rect 800 23056 199200 24136
rect 880 22776 199200 23056
rect 800 21696 199200 22776
rect 880 21416 199200 21696
rect 800 20472 199200 21416
rect 880 20200 199200 20472
rect 880 20192 199120 20200
rect 800 19920 199120 20192
rect 800 19112 199200 19920
rect 880 18832 199200 19112
rect 800 17752 199200 18832
rect 880 17472 199200 17752
rect 800 16528 199200 17472
rect 880 16248 199200 16528
rect 800 15168 199200 16248
rect 880 14888 199200 15168
rect 800 13808 199200 14888
rect 880 13528 199200 13808
rect 800 12584 199200 13528
rect 880 12304 199200 12584
rect 800 11224 199200 12304
rect 880 10944 199200 11224
rect 800 9864 199200 10944
rect 880 9584 199200 9864
rect 800 8640 199200 9584
rect 880 8360 199200 8640
rect 800 7280 199200 8360
rect 880 7000 199200 7280
rect 800 5920 199200 7000
rect 880 5640 199200 5920
rect 800 4696 199200 5640
rect 880 4416 199200 4696
rect 800 3336 199200 4416
rect 880 3056 199200 3336
rect 800 1976 199200 3056
rect 880 1696 199200 1976
rect 800 752 199200 1696
rect 880 579 199200 752
<< metal4 >>
rect 4208 2128 4528 397712
rect 19568 2128 19888 397712
rect 34928 2128 35248 397712
rect 50288 2128 50608 397712
rect 65648 2128 65968 397712
rect 81008 2128 81328 397712
rect 96368 2128 96688 397712
rect 111728 2128 112048 397712
rect 127088 2128 127408 397712
rect 142448 2128 142768 397712
rect 157808 2128 158128 397712
rect 173168 2128 173488 397712
rect 188528 2128 188848 397712
<< obsm4 >>
rect 1347 3435 4128 357509
rect 4608 3435 19488 357509
rect 19968 3435 34848 357509
rect 35328 3435 50208 357509
rect 50688 3435 65568 357509
rect 66048 3435 80901 357509
<< labels >>
rlabel metal3 s 0 174224 800 174344 6 bb_addr0[0]
port 1 nsew signal output
rlabel metal3 s 0 245216 800 245336 6 bb_addr0[10]
port 2 nsew signal output
rlabel metal3 s 0 251744 800 251864 6 bb_addr0[11]
port 3 nsew signal output
rlabel metal3 s 0 258408 800 258528 6 bb_addr0[12]
port 4 nsew signal output
rlabel metal3 s 0 264936 800 265056 6 bb_addr0[13]
port 5 nsew signal output
rlabel metal3 s 0 271464 800 271584 6 bb_addr0[14]
port 6 nsew signal output
rlabel metal3 s 0 278128 800 278248 6 bb_addr0[15]
port 7 nsew signal output
rlabel metal3 s 0 284656 800 284776 6 bb_addr0[16]
port 8 nsew signal output
rlabel metal3 s 0 291320 800 291440 6 bb_addr0[17]
port 9 nsew signal output
rlabel metal3 s 0 297848 800 297968 6 bb_addr0[18]
port 10 nsew signal output
rlabel metal3 s 0 304376 800 304496 6 bb_addr0[19]
port 11 nsew signal output
rlabel metal3 s 0 182112 800 182232 6 bb_addr0[1]
port 12 nsew signal output
rlabel metal3 s 0 311040 800 311160 6 bb_addr0[20]
port 13 nsew signal output
rlabel metal3 s 0 317568 800 317688 6 bb_addr0[21]
port 14 nsew signal output
rlabel metal3 s 0 324096 800 324216 6 bb_addr0[22]
port 15 nsew signal output
rlabel metal3 s 0 330760 800 330880 6 bb_addr0[23]
port 16 nsew signal output
rlabel metal3 s 0 337288 800 337408 6 bb_addr0[24]
port 17 nsew signal output
rlabel metal3 s 0 343952 800 344072 6 bb_addr0[25]
port 18 nsew signal output
rlabel metal3 s 0 350480 800 350600 6 bb_addr0[26]
port 19 nsew signal output
rlabel metal3 s 0 357008 800 357128 6 bb_addr0[27]
port 20 nsew signal output
rlabel metal3 s 0 363672 800 363792 6 bb_addr0[28]
port 21 nsew signal output
rlabel metal3 s 0 370200 800 370320 6 bb_addr0[29]
port 22 nsew signal output
rlabel metal3 s 0 190000 800 190120 6 bb_addr0[2]
port 23 nsew signal output
rlabel metal3 s 0 376728 800 376848 6 bb_addr0[30]
port 24 nsew signal output
rlabel metal3 s 0 383392 800 383512 6 bb_addr0[31]
port 25 nsew signal output
rlabel metal3 s 0 197888 800 198008 6 bb_addr0[3]
port 26 nsew signal output
rlabel metal3 s 0 205776 800 205896 6 bb_addr0[4]
port 27 nsew signal output
rlabel metal3 s 0 212304 800 212424 6 bb_addr0[5]
port 28 nsew signal output
rlabel metal3 s 0 218832 800 218952 6 bb_addr0[6]
port 29 nsew signal output
rlabel metal3 s 0 225496 800 225616 6 bb_addr0[7]
port 30 nsew signal output
rlabel metal3 s 0 232024 800 232144 6 bb_addr0[8]
port 31 nsew signal output
rlabel metal3 s 0 238688 800 238808 6 bb_addr0[9]
port 32 nsew signal output
rlabel metal3 s 0 175448 800 175568 6 bb_addr1[0]
port 33 nsew signal output
rlabel metal3 s 0 246576 800 246696 6 bb_addr1[10]
port 34 nsew signal output
rlabel metal3 s 0 253104 800 253224 6 bb_addr1[11]
port 35 nsew signal output
rlabel metal3 s 0 259632 800 259752 6 bb_addr1[12]
port 36 nsew signal output
rlabel metal3 s 0 266296 800 266416 6 bb_addr1[13]
port 37 nsew signal output
rlabel metal3 s 0 272824 800 272944 6 bb_addr1[14]
port 38 nsew signal output
rlabel metal3 s 0 279352 800 279472 6 bb_addr1[15]
port 39 nsew signal output
rlabel metal3 s 0 286016 800 286136 6 bb_addr1[16]
port 40 nsew signal output
rlabel metal3 s 0 292544 800 292664 6 bb_addr1[17]
port 41 nsew signal output
rlabel metal3 s 0 299208 800 299328 6 bb_addr1[18]
port 42 nsew signal output
rlabel metal3 s 0 305736 800 305856 6 bb_addr1[19]
port 43 nsew signal output
rlabel metal3 s 0 183336 800 183456 6 bb_addr1[1]
port 44 nsew signal output
rlabel metal3 s 0 312264 800 312384 6 bb_addr1[20]
port 45 nsew signal output
rlabel metal3 s 0 318928 800 319048 6 bb_addr1[21]
port 46 nsew signal output
rlabel metal3 s 0 325456 800 325576 6 bb_addr1[22]
port 47 nsew signal output
rlabel metal3 s 0 331984 800 332104 6 bb_addr1[23]
port 48 nsew signal output
rlabel metal3 s 0 338648 800 338768 6 bb_addr1[24]
port 49 nsew signal output
rlabel metal3 s 0 345176 800 345296 6 bb_addr1[25]
port 50 nsew signal output
rlabel metal3 s 0 351840 800 351960 6 bb_addr1[26]
port 51 nsew signal output
rlabel metal3 s 0 358368 800 358488 6 bb_addr1[27]
port 52 nsew signal output
rlabel metal3 s 0 364896 800 365016 6 bb_addr1[28]
port 53 nsew signal output
rlabel metal3 s 0 371560 800 371680 6 bb_addr1[29]
port 54 nsew signal output
rlabel metal3 s 0 191224 800 191344 6 bb_addr1[2]
port 55 nsew signal output
rlabel metal3 s 0 378088 800 378208 6 bb_addr1[30]
port 56 nsew signal output
rlabel metal3 s 0 384616 800 384736 6 bb_addr1[31]
port 57 nsew signal output
rlabel metal3 s 0 199112 800 199232 6 bb_addr1[3]
port 58 nsew signal output
rlabel metal3 s 0 207000 800 207120 6 bb_addr1[4]
port 59 nsew signal output
rlabel metal3 s 0 213664 800 213784 6 bb_addr1[5]
port 60 nsew signal output
rlabel metal3 s 0 220192 800 220312 6 bb_addr1[6]
port 61 nsew signal output
rlabel metal3 s 0 226720 800 226840 6 bb_addr1[7]
port 62 nsew signal output
rlabel metal3 s 0 233384 800 233504 6 bb_addr1[8]
port 63 nsew signal output
rlabel metal3 s 0 239912 800 240032 6 bb_addr1[9]
port 64 nsew signal output
rlabel metal3 s 0 170144 800 170264 6 bb_csb0
port 65 nsew signal output
rlabel metal3 s 0 171504 800 171624 6 bb_csb1
port 66 nsew signal output
rlabel metal3 s 0 176808 800 176928 6 bb_din0[0]
port 67 nsew signal output
rlabel metal3 s 0 247800 800 247920 6 bb_din0[10]
port 68 nsew signal output
rlabel metal3 s 0 254464 800 254584 6 bb_din0[11]
port 69 nsew signal output
rlabel metal3 s 0 260992 800 261112 6 bb_din0[12]
port 70 nsew signal output
rlabel metal3 s 0 267520 800 267640 6 bb_din0[13]
port 71 nsew signal output
rlabel metal3 s 0 274184 800 274304 6 bb_din0[14]
port 72 nsew signal output
rlabel metal3 s 0 280712 800 280832 6 bb_din0[15]
port 73 nsew signal output
rlabel metal3 s 0 287376 800 287496 6 bb_din0[16]
port 74 nsew signal output
rlabel metal3 s 0 293904 800 294024 6 bb_din0[17]
port 75 nsew signal output
rlabel metal3 s 0 300432 800 300552 6 bb_din0[18]
port 76 nsew signal output
rlabel metal3 s 0 307096 800 307216 6 bb_din0[19]
port 77 nsew signal output
rlabel metal3 s 0 184696 800 184816 6 bb_din0[1]
port 78 nsew signal output
rlabel metal3 s 0 313624 800 313744 6 bb_din0[20]
port 79 nsew signal output
rlabel metal3 s 0 320152 800 320272 6 bb_din0[21]
port 80 nsew signal output
rlabel metal3 s 0 326816 800 326936 6 bb_din0[22]
port 81 nsew signal output
rlabel metal3 s 0 333344 800 333464 6 bb_din0[23]
port 82 nsew signal output
rlabel metal3 s 0 339872 800 339992 6 bb_din0[24]
port 83 nsew signal output
rlabel metal3 s 0 346536 800 346656 6 bb_din0[25]
port 84 nsew signal output
rlabel metal3 s 0 353064 800 353184 6 bb_din0[26]
port 85 nsew signal output
rlabel metal3 s 0 359728 800 359848 6 bb_din0[27]
port 86 nsew signal output
rlabel metal3 s 0 366256 800 366376 6 bb_din0[28]
port 87 nsew signal output
rlabel metal3 s 0 372784 800 372904 6 bb_din0[29]
port 88 nsew signal output
rlabel metal3 s 0 192584 800 192704 6 bb_din0[2]
port 89 nsew signal output
rlabel metal3 s 0 379448 800 379568 6 bb_din0[30]
port 90 nsew signal output
rlabel metal3 s 0 385976 800 386096 6 bb_din0[31]
port 91 nsew signal output
rlabel metal3 s 0 200472 800 200592 6 bb_din0[3]
port 92 nsew signal output
rlabel metal3 s 0 208360 800 208480 6 bb_din0[4]
port 93 nsew signal output
rlabel metal3 s 0 214888 800 215008 6 bb_din0[5]
port 94 nsew signal output
rlabel metal3 s 0 221552 800 221672 6 bb_din0[6]
port 95 nsew signal output
rlabel metal3 s 0 228080 800 228200 6 bb_din0[7]
port 96 nsew signal output
rlabel metal3 s 0 234744 800 234864 6 bb_din0[8]
port 97 nsew signal output
rlabel metal3 s 0 241272 800 241392 6 bb_din0[9]
port 98 nsew signal output
rlabel metal3 s 0 178168 800 178288 6 bb_dout0[0]
port 99 nsew signal input
rlabel metal3 s 0 249160 800 249280 6 bb_dout0[10]
port 100 nsew signal input
rlabel metal3 s 0 255688 800 255808 6 bb_dout0[11]
port 101 nsew signal input
rlabel metal3 s 0 262352 800 262472 6 bb_dout0[12]
port 102 nsew signal input
rlabel metal3 s 0 268880 800 269000 6 bb_dout0[13]
port 103 nsew signal input
rlabel metal3 s 0 275408 800 275528 6 bb_dout0[14]
port 104 nsew signal input
rlabel metal3 s 0 282072 800 282192 6 bb_dout0[15]
port 105 nsew signal input
rlabel metal3 s 0 288600 800 288720 6 bb_dout0[16]
port 106 nsew signal input
rlabel metal3 s 0 295264 800 295384 6 bb_dout0[17]
port 107 nsew signal input
rlabel metal3 s 0 301792 800 301912 6 bb_dout0[18]
port 108 nsew signal input
rlabel metal3 s 0 308320 800 308440 6 bb_dout0[19]
port 109 nsew signal input
rlabel metal3 s 0 186056 800 186176 6 bb_dout0[1]
port 110 nsew signal input
rlabel metal3 s 0 314984 800 315104 6 bb_dout0[20]
port 111 nsew signal input
rlabel metal3 s 0 321512 800 321632 6 bb_dout0[21]
port 112 nsew signal input
rlabel metal3 s 0 328040 800 328160 6 bb_dout0[22]
port 113 nsew signal input
rlabel metal3 s 0 334704 800 334824 6 bb_dout0[23]
port 114 nsew signal input
rlabel metal3 s 0 341232 800 341352 6 bb_dout0[24]
port 115 nsew signal input
rlabel metal3 s 0 347896 800 348016 6 bb_dout0[25]
port 116 nsew signal input
rlabel metal3 s 0 354424 800 354544 6 bb_dout0[26]
port 117 nsew signal input
rlabel metal3 s 0 360952 800 361072 6 bb_dout0[27]
port 118 nsew signal input
rlabel metal3 s 0 367616 800 367736 6 bb_dout0[28]
port 119 nsew signal input
rlabel metal3 s 0 374144 800 374264 6 bb_dout0[29]
port 120 nsew signal input
rlabel metal3 s 0 193944 800 194064 6 bb_dout0[2]
port 121 nsew signal input
rlabel metal3 s 0 380672 800 380792 6 bb_dout0[30]
port 122 nsew signal input
rlabel metal3 s 0 387336 800 387456 6 bb_dout0[31]
port 123 nsew signal input
rlabel metal3 s 0 201832 800 201952 6 bb_dout0[3]
port 124 nsew signal input
rlabel metal3 s 0 209720 800 209840 6 bb_dout0[4]
port 125 nsew signal input
rlabel metal3 s 0 216248 800 216368 6 bb_dout0[5]
port 126 nsew signal input
rlabel metal3 s 0 222776 800 222896 6 bb_dout0[6]
port 127 nsew signal input
rlabel metal3 s 0 229440 800 229560 6 bb_dout0[7]
port 128 nsew signal input
rlabel metal3 s 0 235968 800 236088 6 bb_dout0[8]
port 129 nsew signal input
rlabel metal3 s 0 242632 800 242752 6 bb_dout0[9]
port 130 nsew signal input
rlabel metal3 s 0 179392 800 179512 6 bb_dout1[0]
port 131 nsew signal input
rlabel metal3 s 0 250520 800 250640 6 bb_dout1[10]
port 132 nsew signal input
rlabel metal3 s 0 257048 800 257168 6 bb_dout1[11]
port 133 nsew signal input
rlabel metal3 s 0 263576 800 263696 6 bb_dout1[12]
port 134 nsew signal input
rlabel metal3 s 0 270240 800 270360 6 bb_dout1[13]
port 135 nsew signal input
rlabel metal3 s 0 276768 800 276888 6 bb_dout1[14]
port 136 nsew signal input
rlabel metal3 s 0 283296 800 283416 6 bb_dout1[15]
port 137 nsew signal input
rlabel metal3 s 0 289960 800 290080 6 bb_dout1[16]
port 138 nsew signal input
rlabel metal3 s 0 296488 800 296608 6 bb_dout1[17]
port 139 nsew signal input
rlabel metal3 s 0 303152 800 303272 6 bb_dout1[18]
port 140 nsew signal input
rlabel metal3 s 0 309680 800 309800 6 bb_dout1[19]
port 141 nsew signal input
rlabel metal3 s 0 187280 800 187400 6 bb_dout1[1]
port 142 nsew signal input
rlabel metal3 s 0 316208 800 316328 6 bb_dout1[20]
port 143 nsew signal input
rlabel metal3 s 0 322872 800 322992 6 bb_dout1[21]
port 144 nsew signal input
rlabel metal3 s 0 329400 800 329520 6 bb_dout1[22]
port 145 nsew signal input
rlabel metal3 s 0 335928 800 336048 6 bb_dout1[23]
port 146 nsew signal input
rlabel metal3 s 0 342592 800 342712 6 bb_dout1[24]
port 147 nsew signal input
rlabel metal3 s 0 349120 800 349240 6 bb_dout1[25]
port 148 nsew signal input
rlabel metal3 s 0 355784 800 355904 6 bb_dout1[26]
port 149 nsew signal input
rlabel metal3 s 0 362312 800 362432 6 bb_dout1[27]
port 150 nsew signal input
rlabel metal3 s 0 368840 800 368960 6 bb_dout1[28]
port 151 nsew signal input
rlabel metal3 s 0 375504 800 375624 6 bb_dout1[29]
port 152 nsew signal input
rlabel metal3 s 0 195168 800 195288 6 bb_dout1[2]
port 153 nsew signal input
rlabel metal3 s 0 382032 800 382152 6 bb_dout1[30]
port 154 nsew signal input
rlabel metal3 s 0 388560 800 388680 6 bb_dout1[31]
port 155 nsew signal input
rlabel metal3 s 0 203056 800 203176 6 bb_dout1[3]
port 156 nsew signal input
rlabel metal3 s 0 210944 800 211064 6 bb_dout1[4]
port 157 nsew signal input
rlabel metal3 s 0 217608 800 217728 6 bb_dout1[5]
port 158 nsew signal input
rlabel metal3 s 0 224136 800 224256 6 bb_dout1[6]
port 159 nsew signal input
rlabel metal3 s 0 230800 800 230920 6 bb_dout1[7]
port 160 nsew signal input
rlabel metal3 s 0 237328 800 237448 6 bb_dout1[8]
port 161 nsew signal input
rlabel metal3 s 0 243856 800 243976 6 bb_dout1[9]
port 162 nsew signal input
rlabel metal3 s 0 172864 800 172984 6 bb_web0
port 163 nsew signal output
rlabel metal3 s 0 180752 800 180872 6 bb_wmask0[0]
port 164 nsew signal output
rlabel metal3 s 0 188640 800 188760 6 bb_wmask0[1]
port 165 nsew signal output
rlabel metal3 s 0 196528 800 196648 6 bb_wmask0[2]
port 166 nsew signal output
rlabel metal3 s 0 204416 800 204536 6 bb_wmask0[3]
port 167 nsew signal output
rlabel metal2 s 69110 0 69166 800 6 bbb_buy_gecerli_g_w
port 168 nsew signal output
rlabel metal2 s 84566 0 84622 800 6 bbb_buy_ps_g_w[0]
port 169 nsew signal output
rlabel metal3 s 199200 59984 200000 60104 6 bbb_buy_ps_g_w[10]
port 170 nsew signal output
rlabel metal2 s 161478 0 161534 800 6 bbb_buy_ps_g_w[11]
port 171 nsew signal output
rlabel metal2 s 176842 0 176898 800 6 bbb_buy_ps_g_w[12]
port 172 nsew signal output
rlabel metal3 s 0 392504 800 392624 6 bbb_buy_ps_g_w[13]
port 173 nsew signal output
rlabel metal3 s 199200 99968 200000 100088 6 bbb_buy_ps_g_w[14]
port 174 nsew signal output
rlabel metal3 s 199200 139952 200000 140072 6 bbb_buy_ps_g_w[15]
port 175 nsew signal output
rlabel metal3 s 0 393864 800 393984 6 bbb_buy_ps_g_w[16]
port 176 nsew signal output
rlabel metal3 s 199200 179936 200000 180056 6 bbb_buy_ps_g_w[17]
port 177 nsew signal output
rlabel metal3 s 0 395224 800 395344 6 bbb_buy_ps_g_w[18]
port 178 nsew signal output
rlabel metal2 s 192206 0 192262 800 6 bbb_buy_ps_g_w[19]
port 179 nsew signal output
rlabel metal3 s 199200 20000 200000 20120 6 bbb_buy_ps_g_w[1]
port 180 nsew signal output
rlabel metal3 s 199200 219920 200000 220040 6 bbb_buy_ps_g_w[20]
port 181 nsew signal output
rlabel metal3 s 199200 259904 200000 260024 6 bbb_buy_ps_g_w[21]
port 182 nsew signal output
rlabel metal2 s 83278 399200 83334 400000 6 bbb_buy_ps_g_w[22]
port 183 nsew signal output
rlabel metal3 s 0 396448 800 396568 6 bbb_buy_ps_g_w[23]
port 184 nsew signal output
rlabel metal3 s 0 397808 800 397928 6 bbb_buy_ps_g_w[24]
port 185 nsew signal output
rlabel metal3 s 199200 299888 200000 300008 6 bbb_buy_ps_g_w[25]
port 186 nsew signal output
rlabel metal2 s 116674 399200 116730 400000 6 bbb_buy_ps_g_w[26]
port 187 nsew signal output
rlabel metal3 s 0 399168 800 399288 6 bbb_buy_ps_g_w[27]
port 188 nsew signal output
rlabel metal2 s 149978 399200 150034 400000 6 bbb_buy_ps_g_w[28]
port 189 nsew signal output
rlabel metal3 s 199200 339872 200000 339992 6 bbb_buy_ps_g_w[29]
port 190 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 bbb_buy_ps_g_w[2]
port 191 nsew signal output
rlabel metal2 s 183282 399200 183338 400000 6 bbb_buy_ps_g_w[30]
port 192 nsew signal output
rlabel metal3 s 199200 379856 200000 379976 6 bbb_buy_ps_g_w[31]
port 193 nsew signal output
rlabel metal2 s 16670 399200 16726 400000 6 bbb_buy_ps_g_w[3]
port 194 nsew signal output
rlabel metal2 s 49974 399200 50030 400000 6 bbb_buy_ps_g_w[4]
port 195 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 bbb_buy_ps_g_w[5]
port 196 nsew signal output
rlabel metal3 s 0 389920 800 390040 6 bbb_buy_ps_g_w[6]
port 197 nsew signal output
rlabel metal3 s 0 391280 800 391400 6 bbb_buy_ps_g_w[7]
port 198 nsew signal output
rlabel metal2 s 130658 0 130714 800 6 bbb_buy_ps_g_w[8]
port 199 nsew signal output
rlabel metal2 s 146114 0 146170 800 6 bbb_buy_ps_g_w[9]
port 200 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 clk_g
port 201 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 rst_g
port 202 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 rx
port 203 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 tx
port 204 nsew signal output
rlabel metal3 s 0 4496 800 4616 6 vb_addr0[0]
port 205 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 vb_addr0[10]
port 206 nsew signal output
rlabel metal3 s 0 82016 800 82136 6 vb_addr0[11]
port 207 nsew signal output
rlabel metal3 s 0 88680 800 88800 6 vb_addr0[12]
port 208 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 vb_addr0[1]
port 209 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 vb_addr0[2]
port 210 nsew signal output
rlabel metal3 s 0 28160 800 28280 6 vb_addr0[3]
port 211 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 vb_addr0[4]
port 212 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 vb_addr0[5]
port 213 nsew signal output
rlabel metal3 s 0 49104 800 49224 6 vb_addr0[6]
port 214 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 vb_addr0[7]
port 215 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 vb_addr0[8]
port 216 nsew signal output
rlabel metal3 s 0 68960 800 69080 6 vb_addr0[9]
port 217 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 vb_addr1[0]
port 218 nsew signal output
rlabel metal3 s 0 76848 800 76968 6 vb_addr1[10]
port 219 nsew signal output
rlabel metal3 s 0 83376 800 83496 6 vb_addr1[11]
port 220 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 vb_addr1[12]
port 221 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 vb_addr1[1]
port 222 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 vb_addr1[2]
port 223 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 vb_addr1[3]
port 224 nsew signal output
rlabel metal3 s 0 37272 800 37392 6 vb_addr1[4]
port 225 nsew signal output
rlabel metal3 s 0 43936 800 44056 6 vb_addr1[5]
port 226 nsew signal output
rlabel metal3 s 0 50464 800 50584 6 vb_addr1[6]
port 227 nsew signal output
rlabel metal3 s 0 56992 800 57112 6 vb_addr1[7]
port 228 nsew signal output
rlabel metal3 s 0 63656 800 63776 6 vb_addr1[8]
port 229 nsew signal output
rlabel metal3 s 0 70184 800 70304 6 vb_addr1[9]
port 230 nsew signal output
rlabel metal3 s 0 552 800 672 6 vb_csb0
port 231 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 vb_csb1
port 232 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 vb_din0[0]
port 233 nsew signal output
rlabel metal3 s 0 78072 800 78192 6 vb_din0[10]
port 234 nsew signal output
rlabel metal3 s 0 84736 800 84856 6 vb_din0[11]
port 235 nsew signal output
rlabel metal3 s 0 91264 800 91384 6 vb_din0[12]
port 236 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 vb_din0[13]
port 237 nsew signal output
rlabel metal3 s 0 99152 800 99272 6 vb_din0[14]
port 238 nsew signal output
rlabel metal3 s 0 103096 800 103216 6 vb_din0[15]
port 239 nsew signal output
rlabel metal3 s 0 107040 800 107160 6 vb_din0[16]
port 240 nsew signal output
rlabel metal3 s 0 110984 800 111104 6 vb_din0[17]
port 241 nsew signal output
rlabel metal3 s 0 114928 800 115048 6 vb_din0[18]
port 242 nsew signal output
rlabel metal3 s 0 118872 800 118992 6 vb_din0[19]
port 243 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 vb_din0[1]
port 244 nsew signal output
rlabel metal3 s 0 122816 800 122936 6 vb_din0[20]
port 245 nsew signal output
rlabel metal3 s 0 126760 800 126880 6 vb_din0[21]
port 246 nsew signal output
rlabel metal3 s 0 130704 800 130824 6 vb_din0[22]
port 247 nsew signal output
rlabel metal3 s 0 134648 800 134768 6 vb_din0[23]
port 248 nsew signal output
rlabel metal3 s 0 138592 800 138712 6 vb_din0[24]
port 249 nsew signal output
rlabel metal3 s 0 142536 800 142656 6 vb_din0[25]
port 250 nsew signal output
rlabel metal3 s 0 146480 800 146600 6 vb_din0[26]
port 251 nsew signal output
rlabel metal3 s 0 150424 800 150544 6 vb_din0[27]
port 252 nsew signal output
rlabel metal3 s 0 154368 800 154488 6 vb_din0[28]
port 253 nsew signal output
rlabel metal3 s 0 158312 800 158432 6 vb_din0[29]
port 254 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 vb_din0[2]
port 255 nsew signal output
rlabel metal3 s 0 162256 800 162376 6 vb_din0[30]
port 256 nsew signal output
rlabel metal3 s 0 166200 800 166320 6 vb_din0[31]
port 257 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 vb_din0[3]
port 258 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 vb_din0[4]
port 259 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 vb_din0[5]
port 260 nsew signal output
rlabel metal3 s 0 51824 800 51944 6 vb_din0[6]
port 261 nsew signal output
rlabel metal3 s 0 58352 800 58472 6 vb_din0[7]
port 262 nsew signal output
rlabel metal3 s 0 65016 800 65136 6 vb_din0[8]
port 263 nsew signal output
rlabel metal3 s 0 71544 800 71664 6 vb_din0[9]
port 264 nsew signal output
rlabel metal3 s 0 8440 800 8560 6 vb_dout0[0]
port 265 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 vb_dout0[10]
port 266 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 vb_dout0[11]
port 267 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 vb_dout0[12]
port 268 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 vb_dout0[13]
port 269 nsew signal input
rlabel metal3 s 0 100512 800 100632 6 vb_dout0[14]
port 270 nsew signal input
rlabel metal3 s 0 104456 800 104576 6 vb_dout0[15]
port 271 nsew signal input
rlabel metal3 s 0 108400 800 108520 6 vb_dout0[16]
port 272 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 vb_dout0[17]
port 273 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 vb_dout0[18]
port 274 nsew signal input
rlabel metal3 s 0 120232 800 120352 6 vb_dout0[19]
port 275 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 vb_dout0[1]
port 276 nsew signal input
rlabel metal3 s 0 124176 800 124296 6 vb_dout0[20]
port 277 nsew signal input
rlabel metal3 s 0 128120 800 128240 6 vb_dout0[21]
port 278 nsew signal input
rlabel metal3 s 0 132064 800 132184 6 vb_dout0[22]
port 279 nsew signal input
rlabel metal3 s 0 136008 800 136128 6 vb_dout0[23]
port 280 nsew signal input
rlabel metal3 s 0 139952 800 140072 6 vb_dout0[24]
port 281 nsew signal input
rlabel metal3 s 0 143896 800 144016 6 vb_dout0[25]
port 282 nsew signal input
rlabel metal3 s 0 147840 800 147960 6 vb_dout0[26]
port 283 nsew signal input
rlabel metal3 s 0 151784 800 151904 6 vb_dout0[27]
port 284 nsew signal input
rlabel metal3 s 0 155728 800 155848 6 vb_dout0[28]
port 285 nsew signal input
rlabel metal3 s 0 159672 800 159792 6 vb_dout0[29]
port 286 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 vb_dout0[2]
port 287 nsew signal input
rlabel metal3 s 0 163616 800 163736 6 vb_dout0[30]
port 288 nsew signal input
rlabel metal3 s 0 167560 800 167680 6 vb_dout0[31]
port 289 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 vb_dout0[3]
port 290 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 vb_dout0[4]
port 291 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 vb_dout0[5]
port 292 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 vb_dout0[6]
port 293 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 vb_dout0[7]
port 294 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 vb_dout0[8]
port 295 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 vb_dout0[9]
port 296 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 vb_dout1[0]
port 297 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 vb_dout1[10]
port 298 nsew signal input
rlabel metal3 s 0 87320 800 87440 6 vb_dout1[11]
port 299 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 vb_dout1[12]
port 300 nsew signal input
rlabel metal3 s 0 97792 800 97912 6 vb_dout1[13]
port 301 nsew signal input
rlabel metal3 s 0 101736 800 101856 6 vb_dout1[14]
port 302 nsew signal input
rlabel metal3 s 0 105680 800 105800 6 vb_dout1[15]
port 303 nsew signal input
rlabel metal3 s 0 109624 800 109744 6 vb_dout1[16]
port 304 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 vb_dout1[17]
port 305 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 vb_dout1[18]
port 306 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 vb_dout1[19]
port 307 nsew signal input
rlabel metal3 s 0 17552 800 17672 6 vb_dout1[1]
port 308 nsew signal input
rlabel metal3 s 0 125536 800 125656 6 vb_dout1[20]
port 309 nsew signal input
rlabel metal3 s 0 129480 800 129600 6 vb_dout1[21]
port 310 nsew signal input
rlabel metal3 s 0 133424 800 133544 6 vb_dout1[22]
port 311 nsew signal input
rlabel metal3 s 0 137368 800 137488 6 vb_dout1[23]
port 312 nsew signal input
rlabel metal3 s 0 141312 800 141432 6 vb_dout1[24]
port 313 nsew signal input
rlabel metal3 s 0 145256 800 145376 6 vb_dout1[25]
port 314 nsew signal input
rlabel metal3 s 0 149200 800 149320 6 vb_dout1[26]
port 315 nsew signal input
rlabel metal3 s 0 153144 800 153264 6 vb_dout1[27]
port 316 nsew signal input
rlabel metal3 s 0 157088 800 157208 6 vb_dout1[28]
port 317 nsew signal input
rlabel metal3 s 0 161032 800 161152 6 vb_dout1[29]
port 318 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 vb_dout1[2]
port 319 nsew signal input
rlabel metal3 s 0 164976 800 165096 6 vb_dout1[30]
port 320 nsew signal input
rlabel metal3 s 0 168920 800 169040 6 vb_dout1[31]
port 321 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 vb_dout1[3]
port 322 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 vb_dout1[4]
port 323 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 vb_dout1[5]
port 324 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 vb_dout1[6]
port 325 nsew signal input
rlabel metal3 s 0 61072 800 61192 6 vb_dout1[7]
port 326 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 vb_dout1[8]
port 327 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 vb_dout1[9]
port 328 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 vb_web0
port 329 nsew signal output
rlabel metal3 s 0 11024 800 11144 6 vb_wmask0[0]
port 330 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 vb_wmask0[1]
port 331 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 vb_wmask0[2]
port 332 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 vb_wmask0[3]
port 333 nsew signal output
rlabel metal4 s 4208 2128 4528 397712 6 vccd1
port 334 nsew power input
rlabel metal4 s 34928 2128 35248 397712 6 vccd1
port 334 nsew power input
rlabel metal4 s 65648 2128 65968 397712 6 vccd1
port 334 nsew power input
rlabel metal4 s 96368 2128 96688 397712 6 vccd1
port 334 nsew power input
rlabel metal4 s 127088 2128 127408 397712 6 vccd1
port 334 nsew power input
rlabel metal4 s 157808 2128 158128 397712 6 vccd1
port 334 nsew power input
rlabel metal4 s 188528 2128 188848 397712 6 vccd1
port 334 nsew power input
rlabel metal4 s 19568 2128 19888 397712 6 vssd1
port 335 nsew ground input
rlabel metal4 s 50288 2128 50608 397712 6 vssd1
port 335 nsew ground input
rlabel metal4 s 81008 2128 81328 397712 6 vssd1
port 335 nsew ground input
rlabel metal4 s 111728 2128 112048 397712 6 vssd1
port 335 nsew ground input
rlabel metal4 s 142448 2128 142768 397712 6 vssd1
port 335 nsew ground input
rlabel metal4 s 173168 2128 173488 397712 6 vssd1
port 335 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 200000 400000
string LEFview TRUE
string GDS_FILE /home/kasirga/ismail_cup/ismail-mpw4/caravel_user_project/openlane/c0_system_macro/runs/c0_system_macro/results/finishing/c0_system.gds
string GDS_END 78074794
string GDS_START 1266174
<< end >>

