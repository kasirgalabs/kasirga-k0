// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0
`timescale 1ns / 1ps

module c0_uart_prog(
		input c0_tx,
		output reg c0_rx
	);

	// Program len       : 524
	// # of instructions : 111
	// # of data         : 18

	wire [7:0] program [566:0];

	assign program[0] = 8'd188;
	assign program[1] = 8'd1;
	assign program[2] = 8'd0;
	assign program[3] = 8'd0;
	assign program[4] = 8'd111;
	assign program[5] = 8'd0;
	assign program[6] = 8'd128;
	assign program[7] = 8'd4;
	assign program[8] = 8'd115;
	assign program[9] = 8'd47;
	assign program[10] = 8'd32;
	assign program[11] = 8'd52;
	assign program[12] = 8'd147;
	assign program[13] = 8'd15;
	assign program[14] = 8'd128;
	assign program[15] = 8'd0;
	assign program[16] = 8'd99;
	assign program[17] = 8'd8;
	assign program[18] = 8'd255;
	assign program[19] = 8'd3;
	assign program[20] = 8'd147;
	assign program[21] = 8'd15;
	assign program[22] = 8'd144;
	assign program[23] = 8'd0;
	assign program[24] = 8'd99;
	assign program[25] = 8'd4;
	assign program[26] = 8'd255;
	assign program[27] = 8'd3;
	assign program[28] = 8'd147;
	assign program[29] = 8'd15;
	assign program[30] = 8'd176;
	assign program[31] = 8'd0;
	assign program[32] = 8'd99;
	assign program[33] = 8'd0;
	assign program[34] = 8'd255;
	assign program[35] = 8'd3;
	assign program[36] = 8'd19;
	assign program[37] = 8'd15;
	assign program[38] = 8'd0;
	assign program[39] = 8'd0;
	assign program[40] = 8'd99;
	assign program[41] = 8'd4;
	assign program[42] = 8'd15;
	assign program[43] = 8'd0;
	assign program[44] = 8'd103;
	assign program[45] = 8'd0;
	assign program[46] = 8'd15;
	assign program[47] = 8'd0;
	assign program[48] = 8'd115;
	assign program[49] = 8'd47;
	assign program[50] = 8'd32;
	assign program[51] = 8'd52;
	assign program[52] = 8'd99;
	assign program[53] = 8'd84;
	assign program[54] = 8'd15;
	assign program[55] = 8'd0;
	assign program[56] = 8'd111;
	assign program[57] = 8'd0;
	assign program[58] = 8'd64;
	assign program[59] = 8'd0;
	assign program[60] = 8'd147;
	assign program[61] = 8'd225;
	assign program[62] = 8'd145;
	assign program[63] = 8'd83;
	assign program[64] = 8'd23;
	assign program[65] = 8'd15;
	assign program[66] = 8'd31;
	assign program[67] = 8'd0;
	assign program[68] = 8'd35;
	assign program[69] = 8'd34;
	assign program[70] = 8'd63;
	assign program[71] = 8'd252;
	assign program[72] = 8'd111;
	assign program[73] = 8'd240;
	assign program[74] = 8'd159;
	assign program[75] = 8'd255;
	assign program[76] = 8'd147;
	assign program[77] = 8'd0;
	assign program[78] = 8'd0;
	assign program[79] = 8'd0;
	assign program[80] = 8'd19;
	assign program[81] = 8'd1;
	assign program[82] = 8'd0;
	assign program[83] = 8'd0;
	assign program[84] = 8'd147;
	assign program[85] = 8'd1;
	assign program[86] = 8'd0;
	assign program[87] = 8'd0;
	assign program[88] = 8'd19;
	assign program[89] = 8'd2;
	assign program[90] = 8'd0;
	assign program[91] = 8'd0;
	assign program[92] = 8'd147;
	assign program[93] = 8'd2;
	assign program[94] = 8'd0;
	assign program[95] = 8'd0;
	assign program[96] = 8'd19;
	assign program[97] = 8'd3;
	assign program[98] = 8'd0;
	assign program[99] = 8'd0;
	assign program[100] = 8'd147;
	assign program[101] = 8'd3;
	assign program[102] = 8'd0;
	assign program[103] = 8'd0;
	assign program[104] = 8'd19;
	assign program[105] = 8'd4;
	assign program[106] = 8'd0;
	assign program[107] = 8'd0;
	assign program[108] = 8'd147;
	assign program[109] = 8'd4;
	assign program[110] = 8'd0;
	assign program[111] = 8'd0;
	assign program[112] = 8'd19;
	assign program[113] = 8'd5;
	assign program[114] = 8'd0;
	assign program[115] = 8'd0;
	assign program[116] = 8'd147;
	assign program[117] = 8'd5;
	assign program[118] = 8'd0;
	assign program[119] = 8'd0;
	assign program[120] = 8'd19;
	assign program[121] = 8'd6;
	assign program[122] = 8'd0;
	assign program[123] = 8'd0;
	assign program[124] = 8'd147;
	assign program[125] = 8'd6;
	assign program[126] = 8'd0;
	assign program[127] = 8'd0;
	assign program[128] = 8'd19;
	assign program[129] = 8'd7;
	assign program[130] = 8'd0;
	assign program[131] = 8'd0;
	assign program[132] = 8'd147;
	assign program[133] = 8'd7;
	assign program[134] = 8'd0;
	assign program[135] = 8'd0;
	assign program[136] = 8'd19;
	assign program[137] = 8'd8;
	assign program[138] = 8'd0;
	assign program[139] = 8'd0;
	assign program[140] = 8'd147;
	assign program[141] = 8'd8;
	assign program[142] = 8'd0;
	assign program[143] = 8'd0;
	assign program[144] = 8'd19;
	assign program[145] = 8'd9;
	assign program[146] = 8'd0;
	assign program[147] = 8'd0;
	assign program[148] = 8'd147;
	assign program[149] = 8'd9;
	assign program[150] = 8'd0;
	assign program[151] = 8'd0;
	assign program[152] = 8'd19;
	assign program[153] = 8'd10;
	assign program[154] = 8'd0;
	assign program[155] = 8'd0;
	assign program[156] = 8'd147;
	assign program[157] = 8'd10;
	assign program[158] = 8'd0;
	assign program[159] = 8'd0;
	assign program[160] = 8'd19;
	assign program[161] = 8'd11;
	assign program[162] = 8'd0;
	assign program[163] = 8'd0;
	assign program[164] = 8'd147;
	assign program[165] = 8'd11;
	assign program[166] = 8'd0;
	assign program[167] = 8'd0;
	assign program[168] = 8'd19;
	assign program[169] = 8'd12;
	assign program[170] = 8'd0;
	assign program[171] = 8'd0;
	assign program[172] = 8'd147;
	assign program[173] = 8'd12;
	assign program[174] = 8'd0;
	assign program[175] = 8'd0;
	assign program[176] = 8'd19;
	assign program[177] = 8'd13;
	assign program[178] = 8'd0;
	assign program[179] = 8'd0;
	assign program[180] = 8'd147;
	assign program[181] = 8'd13;
	assign program[182] = 8'd0;
	assign program[183] = 8'd0;
	assign program[184] = 8'd19;
	assign program[185] = 8'd14;
	assign program[186] = 8'd0;
	assign program[187] = 8'd0;
	assign program[188] = 8'd147;
	assign program[189] = 8'd14;
	assign program[190] = 8'd0;
	assign program[191] = 8'd0;
	assign program[192] = 8'd19;
	assign program[193] = 8'd15;
	assign program[194] = 8'd0;
	assign program[195] = 8'd0;
	assign program[196] = 8'd147;
	assign program[197] = 8'd15;
	assign program[198] = 8'd0;
	assign program[199] = 8'd0;
	assign program[200] = 8'd115;
	assign program[201] = 8'd37;
	assign program[202] = 8'd64;
	assign program[203] = 8'd241;
	assign program[204] = 8'd99;
	assign program[205] = 8'd16;
	assign program[206] = 8'd5;
	assign program[207] = 8'd0;
	assign program[208] = 8'd151;
	assign program[209] = 8'd2;
	assign program[210] = 8'd0;
	assign program[211] = 8'd0;
	assign program[212] = 8'd147;
	assign program[213] = 8'd130;
	assign program[214] = 8'd2;
	assign program[215] = 8'd1;
	assign program[216] = 8'd115;
	assign program[217] = 8'd144;
	assign program[218] = 8'd82;
	assign program[219] = 8'd48;
	assign program[220] = 8'd115;
	assign program[221] = 8'd80;
	assign program[222] = 8'd0;
	assign program[223] = 8'd24;
	assign program[224] = 8'd151;
	assign program[225] = 8'd2;
	assign program[226] = 8'd0;
	assign program[227] = 8'd0;
	assign program[228] = 8'd147;
	assign program[229] = 8'd130;
	assign program[230] = 8'd2;
	assign program[231] = 8'd2;
	assign program[232] = 8'd115;
	assign program[233] = 8'd144;
	assign program[234] = 8'd82;
	assign program[235] = 8'd48;
	assign program[236] = 8'd183;
	assign program[237] = 8'd2;
	assign program[238] = 8'd0;
	assign program[239] = 8'd128;
	assign program[240] = 8'd147;
	assign program[241] = 8'd130;
	assign program[242] = 8'd242;
	assign program[243] = 8'd255;
	assign program[244] = 8'd115;
	assign program[245] = 8'd144;
	assign program[246] = 8'd2;
	assign program[247] = 8'd59;
	assign program[248] = 8'd147;
	assign program[249] = 8'd2;
	assign program[250] = 8'd240;
	assign program[251] = 8'd1;
	assign program[252] = 8'd115;
	assign program[253] = 8'd144;
	assign program[254] = 8'd2;
	assign program[255] = 8'd58;
	assign program[256] = 8'd115;
	assign program[257] = 8'd80;
	assign program[258] = 8'd64;
	assign program[259] = 8'd48;
	assign program[260] = 8'd151;
	assign program[261] = 8'd2;
	assign program[262] = 8'd0;
	assign program[263] = 8'd0;
	assign program[264] = 8'd147;
	assign program[265] = 8'd130;
	assign program[266] = 8'd66;
	assign program[267] = 8'd1;
	assign program[268] = 8'd115;
	assign program[269] = 8'd144;
	assign program[270] = 8'd82;
	assign program[271] = 8'd48;
	assign program[272] = 8'd115;
	assign program[273] = 8'd80;
	assign program[274] = 8'd32;
	assign program[275] = 8'd48;
	assign program[276] = 8'd115;
	assign program[277] = 8'd80;
	assign program[278] = 8'd48;
	assign program[279] = 8'd48;
	assign program[280] = 8'd147;
	assign program[281] = 8'd1;
	assign program[282] = 8'd0;
	assign program[283] = 8'd0;
	assign program[284] = 8'd151;
	assign program[285] = 8'd2;
	assign program[286] = 8'd0;
	assign program[287] = 8'd0;
	assign program[288] = 8'd147;
	assign program[289] = 8'd130;
	assign program[290] = 8'd194;
	assign program[291] = 8'd238;
	assign program[292] = 8'd115;
	assign program[293] = 8'd144;
	assign program[294] = 8'd82;
	assign program[295] = 8'd48;
	assign program[296] = 8'd19;
	assign program[297] = 8'd5;
	assign program[298] = 8'd16;
	assign program[299] = 8'd0;
	assign program[300] = 8'd19;
	assign program[301] = 8'd21;
	assign program[302] = 8'd245;
	assign program[303] = 8'd1;
	assign program[304] = 8'd99;
	assign program[305] = 8'd76;
	assign program[306] = 8'd5;
	assign program[307] = 8'd0;
	assign program[308] = 8'd15;
	assign program[309] = 8'd0;
	assign program[310] = 8'd240;
	assign program[311] = 8'd15;
	assign program[312] = 8'd147;
	assign program[313] = 8'd1;
	assign program[314] = 8'd16;
	assign program[315] = 8'd0;
	assign program[316] = 8'd147;
	assign program[317] = 8'd8;
	assign program[318] = 8'd208;
	assign program[319] = 8'd5;
	assign program[320] = 8'd19;
	assign program[321] = 8'd5;
	assign program[322] = 8'd0;
	assign program[323] = 8'd0;
	assign program[324] = 8'd115;
	assign program[325] = 8'd0;
	assign program[326] = 8'd0;
	assign program[327] = 8'd0;
	assign program[328] = 8'd147;
	assign program[329] = 8'd2;
	assign program[330] = 8'd0;
	assign program[331] = 8'd0;
	assign program[332] = 8'd99;
	assign program[333] = 8'd138;
	assign program[334] = 8'd2;
	assign program[335] = 8'd0;
	assign program[336] = 8'd115;
	assign program[337] = 8'd144;
	assign program[338] = 8'd82;
	assign program[339] = 8'd16;
	assign program[340] = 8'd183;
	assign program[341] = 8'd178;
	assign program[342] = 8'd0;
	assign program[343] = 8'd0;
	assign program[344] = 8'd147;
	assign program[345] = 8'd130;
	assign program[346] = 8'd146;
	assign program[347] = 8'd16;
	assign program[348] = 8'd115;
	assign program[349] = 8'd144;
	assign program[350] = 8'd34;
	assign program[351] = 8'd48;
	assign program[352] = 8'd115;
	assign program[353] = 8'd80;
	assign program[354] = 8'd0;
	assign program[355] = 8'd48;
	assign program[356] = 8'd151;
	assign program[357] = 8'd2;
	assign program[358] = 8'd0;
	assign program[359] = 8'd0;
	assign program[360] = 8'd147;
	assign program[361] = 8'd130;
	assign program[362] = 8'd66;
	assign program[363] = 8'd1;
	assign program[364] = 8'd115;
	assign program[365] = 8'd144;
	assign program[366] = 8'd18;
	assign program[367] = 8'd52;
	assign program[368] = 8'd115;
	assign program[369] = 8'd37;
	assign program[370] = 8'd64;
	assign program[371] = 8'd241;
	assign program[372] = 8'd115;
	assign program[373] = 8'd0;
	assign program[374] = 8'd32;
	assign program[375] = 8'd48;
	assign program[376] = 8'd15;
	assign program[377] = 8'd0;
	assign program[378] = 8'd240;
	assign program[379] = 8'd15;
	assign program[380] = 8'd147;
	assign program[381] = 8'd1;
	assign program[382] = 8'd16;
	assign program[383] = 8'd0;
	assign program[384] = 8'd147;
	assign program[385] = 8'd8;
	assign program[386] = 8'd208;
	assign program[387] = 8'd5;
	assign program[388] = 8'd19;
	assign program[389] = 8'd5;
	assign program[390] = 8'd0;
	assign program[391] = 8'd0;
	assign program[392] = 8'd115;
	assign program[393] = 8'd0;
	assign program[394] = 8'd0;
	assign program[395] = 8'd0;
	assign program[396] = 8'd115;
	assign program[397] = 8'd16;
	assign program[398] = 8'd0;
	assign program[399] = 8'd192;
	assign program[400] = 8'd0;
	assign program[401] = 8'd0;
	assign program[402] = 8'd0;
	assign program[403] = 8'd0;
	assign program[404] = 8'd0;
	assign program[405] = 8'd0;
	assign program[406] = 8'd0;
	assign program[407] = 8'd0;
	assign program[408] = 8'd0;
	assign program[409] = 8'd0;
	assign program[410] = 8'd0;
	assign program[411] = 8'd0;
	assign program[412] = 8'd0;
	assign program[413] = 8'd0;
	assign program[414] = 8'd0;
	assign program[415] = 8'd0;
	assign program[416] = 8'd0;
	assign program[417] = 8'd0;
	assign program[418] = 8'd0;
	assign program[419] = 8'd0;
	assign program[420] = 8'd0;
	assign program[421] = 8'd0;
	assign program[422] = 8'd0;
	assign program[423] = 8'd0;
	assign program[424] = 8'd0;
	assign program[425] = 8'd0;
	assign program[426] = 8'd0;
	assign program[427] = 8'd0;
	assign program[428] = 8'd0;
	assign program[429] = 8'd0;
	assign program[430] = 8'd0;
	assign program[431] = 8'd0;
	assign program[432] = 8'd0;
	assign program[433] = 8'd0;
	assign program[434] = 8'd0;
	assign program[435] = 8'd0;
	assign program[436] = 8'd0;
	assign program[437] = 8'd0;
	assign program[438] = 8'd0;
	assign program[439] = 8'd0;
	assign program[440] = 8'd0;
	assign program[441] = 8'd0;
	assign program[442] = 8'd0;
	assign program[443] = 8'd0;
	assign program[444] = 8'd0;
	assign program[445] = 8'd0;
	assign program[446] = 8'd0;
	assign program[447] = 8'd0;
	assign program[448] = 8'd72;
	assign program[449] = 8'd0;
	assign program[450] = 8'd0;
	assign program[451] = 8'd0;
	assign program[452] = 8'd0;
	assign program[453] = 8'd0;
	assign program[454] = 8'd0;
	assign program[455] = 8'd0;
	assign program[456] = 8'd0;
	assign program[457] = 8'd0;
	assign program[458] = 8'd0;
	assign program[459] = 8'd0;
	assign program[460] = 8'd0;
	assign program[461] = 8'd0;
	assign program[462] = 8'd0;
	assign program[463] = 8'd0;
	assign program[464] = 8'd0;
	assign program[465] = 8'd0;
	assign program[466] = 8'd0;
	assign program[467] = 8'd0;
	assign program[468] = 8'd0;
	assign program[469] = 8'd0;
	assign program[470] = 8'd0;
	assign program[471] = 8'd0;
	assign program[472] = 8'd0;
	assign program[473] = 8'd0;
	assign program[474] = 8'd0;
	assign program[475] = 8'd0;
	assign program[476] = 8'd0;
	assign program[477] = 8'd0;
	assign program[478] = 8'd0;
	assign program[479] = 8'd0;
	assign program[480] = 8'd0;
	assign program[481] = 8'd0;
	assign program[482] = 8'd0;
	assign program[483] = 8'd0;
	assign program[484] = 8'd0;
	assign program[485] = 8'd0;
	assign program[486] = 8'd0;
	assign program[487] = 8'd0;
	assign program[488] = 8'd0;
	assign program[489] = 8'd0;
	assign program[490] = 8'd0;
	assign program[491] = 8'd0;
	assign program[492] = 8'd0;
	assign program[493] = 8'd0;
	assign program[494] = 8'd0;
	assign program[495] = 8'd0;
	assign program[496] = 8'd0;
	assign program[497] = 8'd0;
	assign program[498] = 8'd0;
	assign program[499] = 8'd0;
	assign program[500] = 8'd0;
	assign program[501] = 8'd0;
	assign program[502] = 8'd0;
	assign program[503] = 8'd0;
	assign program[504] = 8'd0;
	assign program[505] = 8'd0;
	assign program[506] = 8'd0;
	assign program[507] = 8'd0;
	assign program[508] = 8'd0;
	assign program[509] = 8'd0;
	assign program[510] = 8'd0;
	assign program[511] = 8'd0;
	assign program[512] = 8'd0;
	assign program[513] = 8'd0;
	assign program[514] = 8'd0;
	assign program[515] = 8'd0;
	assign program[516] = 8'd0;
	assign program[517] = 8'd0;
	assign program[518] = 8'd0;
	assign program[519] = 8'd0;
	assign program[520] = 8'd0;
	assign program[521] = 8'd0;
	assign program[522] = 8'd0;
	assign program[523] = 8'd0;


	parameter BAUD_PERIOD = 340;
	parameter CLK_PERIOD = 20;

	parameter UART_DELAY = BAUD_PERIOD / CLK_PERIOD;


	integer i, j;
	initial begin
		c0_rx = 1'b1;
		#100000;
		for (i = 0 ; i < 524 ; i = i+1) begin
			c0_rx = 1'b0;
			#BAUD_PERIOD;
			for (j = 0 ; j < 8 ; j = j+1) begin
				c0_rx = program[i][j];
				#BAUD_PERIOD;
			end
			c0_rx = 1'b1;
			#BAUD_PERIOD;
			c0_rx = 1'b1;
			#(BAUD_PERIOD*5);
		end
	end

endmodule
